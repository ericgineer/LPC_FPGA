// top_LPC_FPGA.v

// Generated using ACDS version 15.0 145

`timescale 1 ps / 1 ps
module top_LPC_FPGA (
		output wire        algorithm_run_export,                  //        algorithm_run.export
		output wire        avmm_master_control_rm_fixed_location, //  avmm_master_control.rm_fixed_location
		output wire [31:0] avmm_master_control_rm_read_base,      //                     .rm_read_base
		output wire [31:0] avmm_master_control_rm_read_length,    //                     .rm_read_length
		output wire        avmm_master_control_rm_go,             //                     .rm_go
		input  wire        avmm_master_control_rm_done,           //                     .rm_done
		output wire        avmm_master_control_wm_fixed_location, //                     .wm_fixed_location
		output wire [31:0] avmm_master_control_wm_write_base,     //                     .wm_write_base
		output wire [31:0] avmm_master_control_wm_write_length,   //                     .wm_write_length
		output wire        avmm_master_control_wm_go,             //                     .wm_go
		input  wire        avmm_master_control_wm_done,           //                     .wm_done
		input  wire        clk_clk,                               //                  clk.clk
		output wire [12:0] memory_mem_a,                          //               memory.mem_a
		output wire [2:0]  memory_mem_ba,                         //                     .mem_ba
		output wire [0:0]  memory_mem_ck,                         //                     .mem_ck
		output wire [0:0]  memory_mem_ck_n,                       //                     .mem_ck_n
		output wire [0:0]  memory_mem_cke,                        //                     .mem_cke
		output wire [0:0]  memory_mem_cs_n,                       //                     .mem_cs_n
		output wire [1:0]  memory_mem_dm,                         //                     .mem_dm
		output wire [0:0]  memory_mem_ras_n,                      //                     .mem_ras_n
		output wire [0:0]  memory_mem_cas_n,                      //                     .mem_cas_n
		output wire [0:0]  memory_mem_we_n,                       //                     .mem_we_n
		output wire        memory_mem_reset_n,                    //                     .mem_reset_n
		inout  wire [15:0] memory_mem_dq,                         //                     .mem_dq
		inout  wire [1:0]  memory_mem_dqs,                        //                     .mem_dqs
		inout  wire [1:0]  memory_mem_dqs_n,                      //                     .mem_dqs_n
		output wire [0:0]  memory_mem_odt,                        //                     .mem_odt
		input  wire        oct_rzqin,                             //                  oct.rzqin
		input  wire        read_master_control_fixed_location,    //  read_master_control.fixed_location
		input  wire [31:0] read_master_control_read_base,         //                     .read_base
		input  wire [31:0] read_master_control_read_length,       //                     .read_length
		input  wire        read_master_control_go,                //                     .go
		output wire        read_master_control_done,              //                     .done
		output wire        read_master_control_early_done,        //                     .early_done
		input  wire        read_master_stream_read_buffer,        //   read_master_stream.read_buffer
		output wire [15:0] read_master_stream_buffer_output_data, //                     .buffer_output_data
		output wire        read_master_stream_data_available,     //                     .data_available
		output wire        status_local_init_done,                //               status.local_init_done
		output wire        status_local_cal_success,              //                     .local_cal_success
		output wire        status_local_cal_fail,                 //                     .local_cal_fail
		input  wire        write_master_control_fixed_location,   // write_master_control.fixed_location
		input  wire [31:0] write_master_control_write_base,       //                     .write_base
		input  wire [31:0] write_master_control_write_length,     //                     .write_length
		input  wire        write_master_control_go,               //                     .go
		output wire        write_master_control_done,             //                     .done
		input  wire        write_master_stream_write_buffer,      //  write_master_stream.write_buffer
		input  wire [15:0] write_master_stream_buffer_input_data, //                     .buffer_input_data
		output wire        write_master_stream_buffer_full        //                     .buffer_full
	);

	wire         clk_divide_8k_0_clock_out_clk;                                             // clk_divide_8k_0:clk_out -> [AlgorithmRun:clk, DDR3_interface:mp_cmd_clk_0_clk, DDR3_interface:mp_cmd_clk_1_clk, DDR3_interface:mp_cmd_clk_2_clk, DDR3_interface:mp_rfifo_clk_0_clk, DDR3_interface:mp_rfifo_clk_1_clk, DDR3_interface:mp_rfifo_clk_2_clk, DDR3_interface:mp_wfifo_clk_0_clk, DDR3_interface:mp_wfifo_clk_1_clk, DDR3_interface:mp_wfifo_clk_2_clk, JTAG_master:clk_clk, avmm_master_interface_0:clk, mm_interconnect_0:clk_divide_8k_0_clock_out_clk, mm_interconnect_1:clk_divide_8k_0_clock_out_clk, mm_interconnect_2:clk_divide_8k_0_clock_out_clk, read_master:clk, rst_controller:clk, write_master:clk]
	wire         jtag_master_master_reset_reset;                                            // JTAG_master:master_reset_reset -> [DDR3_interface:global_reset_n, DDR3_interface:mp_cmd_reset_n_0_reset_n, DDR3_interface:mp_cmd_reset_n_1_reset_n, DDR3_interface:mp_cmd_reset_n_2_reset_n, DDR3_interface:mp_rfifo_reset_n_0_reset_n, DDR3_interface:mp_rfifo_reset_n_1_reset_n, DDR3_interface:mp_rfifo_reset_n_2_reset_n, DDR3_interface:mp_wfifo_reset_n_0_reset_n, DDR3_interface:mp_wfifo_reset_n_1_reset_n, DDR3_interface:mp_wfifo_reset_n_2_reset_n, DDR3_interface:soft_reset_n, JTAG_master:clk_reset_reset, rst_controller:reset_in0, rst_controller_001:reset_in0]
	wire  [15:0] read_master_avalon_master_readdata;                                        // mm_interconnect_0:read_master_avalon_master_readdata -> read_master:master_readdata
	wire         read_master_avalon_master_waitrequest;                                     // mm_interconnect_0:read_master_avalon_master_waitrequest -> read_master:master_waitrequest
	wire  [31:0] read_master_avalon_master_address;                                         // read_master:master_address -> mm_interconnect_0:read_master_avalon_master_address
	wire         read_master_avalon_master_read;                                            // read_master:master_read -> mm_interconnect_0:read_master_avalon_master_read
	wire   [1:0] read_master_avalon_master_byteenable;                                      // read_master:master_byteenable -> mm_interconnect_0:read_master_avalon_master_byteenable
	wire         read_master_avalon_master_readdatavalid;                                   // mm_interconnect_0:read_master_avalon_master_readdatavalid -> read_master:master_readdatavalid
	wire   [2:0] read_master_avalon_master_burstcount;                                      // read_master:master_burstcount -> mm_interconnect_0:read_master_avalon_master_burstcount
	wire         mm_interconnect_0_ddr3_interface_avl_1_beginbursttransfer;                 // mm_interconnect_0:DDR3_interface_avl_1_beginbursttransfer -> DDR3_interface:avl_burstbegin_1
	wire  [31:0] mm_interconnect_0_ddr3_interface_avl_1_readdata;                           // DDR3_interface:avl_rdata_1 -> mm_interconnect_0:DDR3_interface_avl_1_readdata
	wire         mm_interconnect_0_ddr3_interface_avl_1_waitrequest;                        // DDR3_interface:avl_ready_1 -> mm_interconnect_0:DDR3_interface_avl_1_waitrequest
	wire  [24:0] mm_interconnect_0_ddr3_interface_avl_1_address;                            // mm_interconnect_0:DDR3_interface_avl_1_address -> DDR3_interface:avl_addr_1
	wire         mm_interconnect_0_ddr3_interface_avl_1_read;                               // mm_interconnect_0:DDR3_interface_avl_1_read -> DDR3_interface:avl_read_req_1
	wire   [3:0] mm_interconnect_0_ddr3_interface_avl_1_byteenable;                         // mm_interconnect_0:DDR3_interface_avl_1_byteenable -> DDR3_interface:avl_be_1
	wire         mm_interconnect_0_ddr3_interface_avl_1_readdatavalid;                      // DDR3_interface:avl_rdata_valid_1 -> mm_interconnect_0:DDR3_interface_avl_1_readdatavalid
	wire         mm_interconnect_0_ddr3_interface_avl_1_write;                              // mm_interconnect_0:DDR3_interface_avl_1_write -> DDR3_interface:avl_write_req_1
	wire  [31:0] mm_interconnect_0_ddr3_interface_avl_1_writedata;                          // mm_interconnect_0:DDR3_interface_avl_1_writedata -> DDR3_interface:avl_wdata_1
	wire   [2:0] mm_interconnect_0_ddr3_interface_avl_1_burstcount;                         // mm_interconnect_0:DDR3_interface_avl_1_burstcount -> DDR3_interface:avl_size_1
	wire         write_master_avalon_master_waitrequest;                                    // mm_interconnect_1:write_master_avalon_master_waitrequest -> write_master:master_waitrequest
	wire  [31:0] write_master_avalon_master_address;                                        // write_master:master_address -> mm_interconnect_1:write_master_avalon_master_address
	wire   [1:0] write_master_avalon_master_byteenable;                                     // write_master:master_byteenable -> mm_interconnect_1:write_master_avalon_master_byteenable
	wire         write_master_avalon_master_write;                                          // write_master:master_write -> mm_interconnect_1:write_master_avalon_master_write
	wire  [15:0] write_master_avalon_master_writedata;                                      // write_master:master_writedata -> mm_interconnect_1:write_master_avalon_master_writedata
	wire   [2:0] write_master_avalon_master_burstcount;                                     // write_master:master_burstcount -> mm_interconnect_1:write_master_avalon_master_burstcount
	wire         mm_interconnect_1_ddr3_interface_avl_2_beginbursttransfer;                 // mm_interconnect_1:DDR3_interface_avl_2_beginbursttransfer -> DDR3_interface:avl_burstbegin_2
	wire  [31:0] mm_interconnect_1_ddr3_interface_avl_2_readdata;                           // DDR3_interface:avl_rdata_2 -> mm_interconnect_1:DDR3_interface_avl_2_readdata
	wire         mm_interconnect_1_ddr3_interface_avl_2_waitrequest;                        // DDR3_interface:avl_ready_2 -> mm_interconnect_1:DDR3_interface_avl_2_waitrequest
	wire  [24:0] mm_interconnect_1_ddr3_interface_avl_2_address;                            // mm_interconnect_1:DDR3_interface_avl_2_address -> DDR3_interface:avl_addr_2
	wire         mm_interconnect_1_ddr3_interface_avl_2_read;                               // mm_interconnect_1:DDR3_interface_avl_2_read -> DDR3_interface:avl_read_req_2
	wire   [3:0] mm_interconnect_1_ddr3_interface_avl_2_byteenable;                         // mm_interconnect_1:DDR3_interface_avl_2_byteenable -> DDR3_interface:avl_be_2
	wire         mm_interconnect_1_ddr3_interface_avl_2_readdatavalid;                      // DDR3_interface:avl_rdata_valid_2 -> mm_interconnect_1:DDR3_interface_avl_2_readdatavalid
	wire         mm_interconnect_1_ddr3_interface_avl_2_write;                              // mm_interconnect_1:DDR3_interface_avl_2_write -> DDR3_interface:avl_write_req_2
	wire  [31:0] mm_interconnect_1_ddr3_interface_avl_2_writedata;                          // mm_interconnect_1:DDR3_interface_avl_2_writedata -> DDR3_interface:avl_wdata_2
	wire   [2:0] mm_interconnect_1_ddr3_interface_avl_2_burstcount;                         // mm_interconnect_1:DDR3_interface_avl_2_burstcount -> DDR3_interface:avl_size_2
	wire  [31:0] jtag_master_master_readdata;                                               // mm_interconnect_2:JTAG_master_master_readdata -> JTAG_master:master_readdata
	wire         jtag_master_master_waitrequest;                                            // mm_interconnect_2:JTAG_master_master_waitrequest -> JTAG_master:master_waitrequest
	wire  [31:0] jtag_master_master_address;                                                // JTAG_master:master_address -> mm_interconnect_2:JTAG_master_master_address
	wire         jtag_master_master_read;                                                   // JTAG_master:master_read -> mm_interconnect_2:JTAG_master_master_read
	wire   [3:0] jtag_master_master_byteenable;                                             // JTAG_master:master_byteenable -> mm_interconnect_2:JTAG_master_master_byteenable
	wire         jtag_master_master_readdatavalid;                                          // mm_interconnect_2:JTAG_master_master_readdatavalid -> JTAG_master:master_readdatavalid
	wire         jtag_master_master_write;                                                  // JTAG_master:master_write -> mm_interconnect_2:JTAG_master_master_write
	wire  [31:0] jtag_master_master_writedata;                                              // JTAG_master:master_writedata -> mm_interconnect_2:JTAG_master_master_writedata
	wire         mm_interconnect_2_ddr3_interface_avl_0_beginbursttransfer;                 // mm_interconnect_2:DDR3_interface_avl_0_beginbursttransfer -> DDR3_interface:avl_burstbegin_0
	wire  [31:0] mm_interconnect_2_ddr3_interface_avl_0_readdata;                           // DDR3_interface:avl_rdata_0 -> mm_interconnect_2:DDR3_interface_avl_0_readdata
	wire         mm_interconnect_2_ddr3_interface_avl_0_waitrequest;                        // DDR3_interface:avl_ready_0 -> mm_interconnect_2:DDR3_interface_avl_0_waitrequest
	wire  [24:0] mm_interconnect_2_ddr3_interface_avl_0_address;                            // mm_interconnect_2:DDR3_interface_avl_0_address -> DDR3_interface:avl_addr_0
	wire         mm_interconnect_2_ddr3_interface_avl_0_read;                               // mm_interconnect_2:DDR3_interface_avl_0_read -> DDR3_interface:avl_read_req_0
	wire   [3:0] mm_interconnect_2_ddr3_interface_avl_0_byteenable;                         // mm_interconnect_2:DDR3_interface_avl_0_byteenable -> DDR3_interface:avl_be_0
	wire         mm_interconnect_2_ddr3_interface_avl_0_readdatavalid;                      // DDR3_interface:avl_rdata_valid_0 -> mm_interconnect_2:DDR3_interface_avl_0_readdatavalid
	wire         mm_interconnect_2_ddr3_interface_avl_0_write;                              // mm_interconnect_2:DDR3_interface_avl_0_write -> DDR3_interface:avl_write_req_0
	wire  [31:0] mm_interconnect_2_ddr3_interface_avl_0_writedata;                          // mm_interconnect_2:DDR3_interface_avl_0_writedata -> DDR3_interface:avl_wdata_0
	wire   [2:0] mm_interconnect_2_ddr3_interface_avl_0_burstcount;                         // mm_interconnect_2:DDR3_interface_avl_0_burstcount -> DDR3_interface:avl_size_0
	wire  [31:0] mm_interconnect_2_avmm_master_interface_0_avmm_master_interface_readdata;  // avmm_master_interface_0:readdata -> mm_interconnect_2:avmm_master_interface_0_avmm_master_interface_readdata
	wire   [3:0] mm_interconnect_2_avmm_master_interface_0_avmm_master_interface_address;   // mm_interconnect_2:avmm_master_interface_0_avmm_master_interface_address -> avmm_master_interface_0:address
	wire         mm_interconnect_2_avmm_master_interface_0_avmm_master_interface_read;      // mm_interconnect_2:avmm_master_interface_0_avmm_master_interface_read -> avmm_master_interface_0:read
	wire         mm_interconnect_2_avmm_master_interface_0_avmm_master_interface_write;     // mm_interconnect_2:avmm_master_interface_0_avmm_master_interface_write -> avmm_master_interface_0:write
	wire  [31:0] mm_interconnect_2_avmm_master_interface_0_avmm_master_interface_writedata; // mm_interconnect_2:avmm_master_interface_0_avmm_master_interface_writedata -> avmm_master_interface_0:writedata
	wire         mm_interconnect_2_algorithmrun_s1_chipselect;                              // mm_interconnect_2:AlgorithmRun_s1_chipselect -> AlgorithmRun:chipselect
	wire  [31:0] mm_interconnect_2_algorithmrun_s1_readdata;                                // AlgorithmRun:readdata -> mm_interconnect_2:AlgorithmRun_s1_readdata
	wire   [1:0] mm_interconnect_2_algorithmrun_s1_address;                                 // mm_interconnect_2:AlgorithmRun_s1_address -> AlgorithmRun:address
	wire         mm_interconnect_2_algorithmrun_s1_write;                                   // mm_interconnect_2:AlgorithmRun_s1_write -> AlgorithmRun:write_n
	wire  [31:0] mm_interconnect_2_algorithmrun_s1_writedata;                               // mm_interconnect_2:AlgorithmRun_s1_writedata -> AlgorithmRun:writedata
	wire         rst_controller_reset_out_reset;                                            // rst_controller:reset_out -> [AlgorithmRun:reset_n, avmm_master_interface_0:rst, mm_interconnect_0:DDR3_interface_mp_cmd_reset_n_1_reset_bridge_in_reset_reset, mm_interconnect_0:read_master_clock_reset_reset_reset_bridge_in_reset_reset, mm_interconnect_1:DDR3_interface_mp_cmd_reset_n_2_reset_bridge_in_reset_reset, mm_interconnect_1:write_master_clock_reset_reset_reset_bridge_in_reset_reset, mm_interconnect_2:JTAG_master_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_2:avmm_master_interface_0_reset_reset_bridge_in_reset_reset, read_master:reset, write_master:reset]
	wire         rst_controller_001_reset_out_reset;                                        // rst_controller_001:reset_out -> clk_divide_8k_0:clk_rst

	top_LPC_FPGA_AlgorithmRun algorithmrun (
		.clk        (clk_divide_8k_0_clock_out_clk),                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_2_algorithmrun_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_2_algorithmrun_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_2_algorithmrun_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_2_algorithmrun_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_2_algorithmrun_s1_readdata),   //                    .readdata
		.out_port   (algorithm_run_export)                          // external_connection.export
	);

	top_LPC_FPGA_DDR3_interface ddr3_interface (
		.pll_ref_clk                (clk_clk),                                                   //        pll_ref_clk.clk
		.global_reset_n             (~jtag_master_master_reset_reset),                           //       global_reset.reset_n
		.soft_reset_n               (~jtag_master_master_reset_reset),                           //         soft_reset.reset_n
		.afi_clk                    (),                                                          //            afi_clk.clk
		.afi_half_clk               (),                                                          //       afi_half_clk.clk
		.afi_reset_n                (),                                                          //          afi_reset.reset_n
		.afi_reset_export_n         (),                                                          //   afi_reset_export.reset_n
		.mem_a                      (memory_mem_a),                                              //             memory.mem_a
		.mem_ba                     (memory_mem_ba),                                             //                   .mem_ba
		.mem_ck                     (memory_mem_ck),                                             //                   .mem_ck
		.mem_ck_n                   (memory_mem_ck_n),                                           //                   .mem_ck_n
		.mem_cke                    (memory_mem_cke),                                            //                   .mem_cke
		.mem_cs_n                   (memory_mem_cs_n),                                           //                   .mem_cs_n
		.mem_dm                     (memory_mem_dm),                                             //                   .mem_dm
		.mem_ras_n                  (memory_mem_ras_n),                                          //                   .mem_ras_n
		.mem_cas_n                  (memory_mem_cas_n),                                          //                   .mem_cas_n
		.mem_we_n                   (memory_mem_we_n),                                           //                   .mem_we_n
		.mem_reset_n                (memory_mem_reset_n),                                        //                   .mem_reset_n
		.mem_dq                     (memory_mem_dq),                                             //                   .mem_dq
		.mem_dqs                    (memory_mem_dqs),                                            //                   .mem_dqs
		.mem_dqs_n                  (memory_mem_dqs_n),                                          //                   .mem_dqs_n
		.mem_odt                    (memory_mem_odt),                                            //                   .mem_odt
		.avl_ready_0                (mm_interconnect_2_ddr3_interface_avl_0_waitrequest),        //              avl_0.waitrequest_n
		.avl_burstbegin_0           (mm_interconnect_2_ddr3_interface_avl_0_beginbursttransfer), //                   .beginbursttransfer
		.avl_addr_0                 (mm_interconnect_2_ddr3_interface_avl_0_address),            //                   .address
		.avl_rdata_valid_0          (mm_interconnect_2_ddr3_interface_avl_0_readdatavalid),      //                   .readdatavalid
		.avl_rdata_0                (mm_interconnect_2_ddr3_interface_avl_0_readdata),           //                   .readdata
		.avl_wdata_0                (mm_interconnect_2_ddr3_interface_avl_0_writedata),          //                   .writedata
		.avl_be_0                   (mm_interconnect_2_ddr3_interface_avl_0_byteenable),         //                   .byteenable
		.avl_read_req_0             (mm_interconnect_2_ddr3_interface_avl_0_read),               //                   .read
		.avl_write_req_0            (mm_interconnect_2_ddr3_interface_avl_0_write),              //                   .write
		.avl_size_0                 (mm_interconnect_2_ddr3_interface_avl_0_burstcount),         //                   .burstcount
		.avl_ready_1                (mm_interconnect_0_ddr3_interface_avl_1_waitrequest),        //              avl_1.waitrequest_n
		.avl_burstbegin_1           (mm_interconnect_0_ddr3_interface_avl_1_beginbursttransfer), //                   .beginbursttransfer
		.avl_addr_1                 (mm_interconnect_0_ddr3_interface_avl_1_address),            //                   .address
		.avl_rdata_valid_1          (mm_interconnect_0_ddr3_interface_avl_1_readdatavalid),      //                   .readdatavalid
		.avl_rdata_1                (mm_interconnect_0_ddr3_interface_avl_1_readdata),           //                   .readdata
		.avl_wdata_1                (mm_interconnect_0_ddr3_interface_avl_1_writedata),          //                   .writedata
		.avl_be_1                   (mm_interconnect_0_ddr3_interface_avl_1_byteenable),         //                   .byteenable
		.avl_read_req_1             (mm_interconnect_0_ddr3_interface_avl_1_read),               //                   .read
		.avl_write_req_1            (mm_interconnect_0_ddr3_interface_avl_1_write),              //                   .write
		.avl_size_1                 (mm_interconnect_0_ddr3_interface_avl_1_burstcount),         //                   .burstcount
		.avl_ready_2                (mm_interconnect_1_ddr3_interface_avl_2_waitrequest),        //              avl_2.waitrequest_n
		.avl_burstbegin_2           (mm_interconnect_1_ddr3_interface_avl_2_beginbursttransfer), //                   .beginbursttransfer
		.avl_addr_2                 (mm_interconnect_1_ddr3_interface_avl_2_address),            //                   .address
		.avl_rdata_valid_2          (mm_interconnect_1_ddr3_interface_avl_2_readdatavalid),      //                   .readdatavalid
		.avl_rdata_2                (mm_interconnect_1_ddr3_interface_avl_2_readdata),           //                   .readdata
		.avl_wdata_2                (mm_interconnect_1_ddr3_interface_avl_2_writedata),          //                   .writedata
		.avl_be_2                   (mm_interconnect_1_ddr3_interface_avl_2_byteenable),         //                   .byteenable
		.avl_read_req_2             (mm_interconnect_1_ddr3_interface_avl_2_read),               //                   .read
		.avl_write_req_2            (mm_interconnect_1_ddr3_interface_avl_2_write),              //                   .write
		.avl_size_2                 (mm_interconnect_1_ddr3_interface_avl_2_burstcount),         //                   .burstcount
		.mp_cmd_clk_0_clk           (clk_divide_8k_0_clock_out_clk),                             //       mp_cmd_clk_0.clk
		.mp_cmd_reset_n_0_reset_n   (~jtag_master_master_reset_reset),                           //   mp_cmd_reset_n_0.reset_n
		.mp_cmd_clk_1_clk           (clk_divide_8k_0_clock_out_clk),                             //       mp_cmd_clk_1.clk
		.mp_cmd_reset_n_1_reset_n   (~jtag_master_master_reset_reset),                           //   mp_cmd_reset_n_1.reset_n
		.mp_cmd_clk_2_clk           (clk_divide_8k_0_clock_out_clk),                             //       mp_cmd_clk_2.clk
		.mp_cmd_reset_n_2_reset_n   (~jtag_master_master_reset_reset),                           //   mp_cmd_reset_n_2.reset_n
		.mp_rfifo_clk_0_clk         (clk_divide_8k_0_clock_out_clk),                             //     mp_rfifo_clk_0.clk
		.mp_rfifo_reset_n_0_reset_n (~jtag_master_master_reset_reset),                           // mp_rfifo_reset_n_0.reset_n
		.mp_wfifo_clk_0_clk         (clk_divide_8k_0_clock_out_clk),                             //     mp_wfifo_clk_0.clk
		.mp_wfifo_reset_n_0_reset_n (~jtag_master_master_reset_reset),                           // mp_wfifo_reset_n_0.reset_n
		.mp_rfifo_clk_1_clk         (clk_divide_8k_0_clock_out_clk),                             //     mp_rfifo_clk_1.clk
		.mp_rfifo_reset_n_1_reset_n (~jtag_master_master_reset_reset),                           // mp_rfifo_reset_n_1.reset_n
		.mp_wfifo_clk_1_clk         (clk_divide_8k_0_clock_out_clk),                             //     mp_wfifo_clk_1.clk
		.mp_wfifo_reset_n_1_reset_n (~jtag_master_master_reset_reset),                           // mp_wfifo_reset_n_1.reset_n
		.mp_rfifo_clk_2_clk         (clk_divide_8k_0_clock_out_clk),                             //     mp_rfifo_clk_2.clk
		.mp_rfifo_reset_n_2_reset_n (~jtag_master_master_reset_reset),                           // mp_rfifo_reset_n_2.reset_n
		.mp_wfifo_clk_2_clk         (clk_divide_8k_0_clock_out_clk),                             //     mp_wfifo_clk_2.clk
		.mp_wfifo_reset_n_2_reset_n (~jtag_master_master_reset_reset),                           // mp_wfifo_reset_n_2.reset_n
		.local_init_done            (status_local_init_done),                                    //             status.local_init_done
		.local_cal_success          (status_local_cal_success),                                  //                   .local_cal_success
		.local_cal_fail             (status_local_cal_fail),                                     //                   .local_cal_fail
		.oct_rzqin                  (oct_rzqin),                                                 //                oct.rzqin
		.pll_mem_clk                (),                                                          //        pll_sharing.pll_mem_clk
		.pll_write_clk              (),                                                          //                   .pll_write_clk
		.pll_locked                 (),                                                          //                   .pll_locked
		.pll_write_clk_pre_phy_clk  (),                                                          //                   .pll_write_clk_pre_phy_clk
		.pll_addr_cmd_clk           (),                                                          //                   .pll_addr_cmd_clk
		.pll_avl_clk                (),                                                          //                   .pll_avl_clk
		.pll_config_clk             (),                                                          //                   .pll_config_clk
		.pll_mem_phy_clk            (),                                                          //                   .pll_mem_phy_clk
		.afi_phy_clk                (),                                                          //                   .afi_phy_clk
		.pll_avl_phy_clk            ()                                                           //                   .pll_avl_phy_clk
	);

	top_LPC_FPGA_JTAG_master #(
		.USE_PLI     (0),
		.PLI_PORT    (50000),
		.FIFO_DEPTHS (2)
	) jtag_master (
		.clk_clk              (clk_divide_8k_0_clock_out_clk),    //          clk.clk
		.clk_reset_reset      (jtag_master_master_reset_reset),   //    clk_reset.reset
		.master_address       (jtag_master_master_address),       //       master.address
		.master_readdata      (jtag_master_master_readdata),      //             .readdata
		.master_read          (jtag_master_master_read),          //             .read
		.master_write         (jtag_master_master_write),         //             .write
		.master_writedata     (jtag_master_master_writedata),     //             .writedata
		.master_waitrequest   (jtag_master_master_waitrequest),   //             .waitrequest
		.master_readdatavalid (jtag_master_master_readdatavalid), //             .readdatavalid
		.master_byteenable    (jtag_master_master_byteenable),    //             .byteenable
		.master_reset_reset   (jtag_master_master_reset_reset)    // master_reset.reset
	);

	master_avalon_interface avmm_master_interface_0 (
		.clk                         (clk_divide_8k_0_clock_out_clk),                                             //                 clock.clk
		.address                     (mm_interconnect_2_avmm_master_interface_0_avmm_master_interface_address),   // avmm_master_interface.address
		.write                       (mm_interconnect_2_avmm_master_interface_0_avmm_master_interface_write),     //                      .write
		.read                        (mm_interconnect_2_avmm_master_interface_0_avmm_master_interface_read),      //                      .read
		.writedata                   (mm_interconnect_2_avmm_master_interface_0_avmm_master_interface_writedata), //                      .writedata
		.readdata                    (mm_interconnect_2_avmm_master_interface_0_avmm_master_interface_readdata),  //                      .readdata
		.read_master_fixed_location  (avmm_master_control_rm_fixed_location),                                     //        master_control.rm_fixed_location
		.read_master_read_base       (avmm_master_control_rm_read_base),                                          //                      .rm_read_base
		.read_master_read_length     (avmm_master_control_rm_read_length),                                        //                      .rm_read_length
		.read_master_go              (avmm_master_control_rm_go),                                                 //                      .rm_go
		.read_master_done            (avmm_master_control_rm_done),                                               //                      .rm_done
		.write_master_fixed_location (avmm_master_control_wm_fixed_location),                                     //                      .wm_fixed_location
		.write_master_write_base     (avmm_master_control_wm_write_base),                                         //                      .wm_write_base
		.write_master_write_length   (avmm_master_control_wm_write_length),                                       //                      .wm_write_length
		.write_master_go             (avmm_master_control_wm_go),                                                 //                      .wm_go
		.write_master_done           (avmm_master_control_wm_done),                                               //                      .wm_done
		.rst                         (rst_controller_reset_out_reset)                                             //                 reset.reset
	);

	clk_divide clk_divide_8k_0 (
		.clk         (clk_clk),                            //           clock.clk
		.clk_out     (clk_divide_8k_0_clock_out_clk),      //       clock_out.clk
		.clk_rst     (rst_controller_001_reset_out_reset), //     clock_reset.reset
		.clk_rst_out ()                                    // clock_reset_out.reset
	);

	custom_master #(
		.MASTER_DIRECTION    (0),
		.DATA_WIDTH          (16),
		.ADDRESS_WIDTH       (32),
		.BURST_CAPABLE       (1),
		.MAXIMUM_BURST_COUNT (4),
		.BURST_COUNT_WIDTH   (3),
		.FIFO_DEPTH          (32),
		.FIFO_DEPTH_LOG2     (5),
		.MEMORY_BASED_FIFO   (1)
	) read_master (
		.clk                     (clk_divide_8k_0_clock_out_clk),           //       clock_reset.clk
		.reset                   (rst_controller_reset_out_reset),          // clock_reset_reset.reset
		.master_address          (read_master_avalon_master_address),       //     avalon_master.address
		.master_read             (read_master_avalon_master_read),          //                  .read
		.master_byteenable       (read_master_avalon_master_byteenable),    //                  .byteenable
		.master_readdata         (read_master_avalon_master_readdata),      //                  .readdata
		.master_readdatavalid    (read_master_avalon_master_readdatavalid), //                  .readdatavalid
		.master_burstcount       (read_master_avalon_master_burstcount),    //                  .burstcount
		.master_waitrequest      (read_master_avalon_master_waitrequest),   //                  .waitrequest
		.control_fixed_location  (read_master_control_fixed_location),      //           control.export
		.control_read_base       (read_master_control_read_base),           //                  .export
		.control_read_length     (read_master_control_read_length),         //                  .export
		.control_go              (read_master_control_go),                  //                  .export
		.control_done            (read_master_control_done),                //                  .export
		.control_early_done      (read_master_control_early_done),          //                  .export
		.user_read_buffer        (read_master_stream_read_buffer),          //              user.export
		.user_buffer_output_data (read_master_stream_buffer_output_data),   //                  .export
		.user_data_available     (read_master_stream_data_available),       //                  .export
		.master_write            (),                                        //       (terminated)
		.master_writedata        (),                                        //       (terminated)
		.control_write_base      (32'b00000000000000000000000000000000),    //       (terminated)
		.control_write_length    (32'b00000000000000000000000000000000),    //       (terminated)
		.user_write_buffer       (1'b0),                                    //       (terminated)
		.user_buffer_input_data  (16'b0000000000000000),                    //       (terminated)
		.user_buffer_full        ()                                         //       (terminated)
	);

	custom_master #(
		.MASTER_DIRECTION    (1),
		.DATA_WIDTH          (16),
		.ADDRESS_WIDTH       (32),
		.BURST_CAPABLE       (1),
		.MAXIMUM_BURST_COUNT (4),
		.BURST_COUNT_WIDTH   (3),
		.FIFO_DEPTH          (32),
		.FIFO_DEPTH_LOG2     (5),
		.MEMORY_BASED_FIFO   (1)
	) write_master (
		.clk                     (clk_divide_8k_0_clock_out_clk),          //       clock_reset.clk
		.reset                   (rst_controller_reset_out_reset),         // clock_reset_reset.reset
		.master_address          (write_master_avalon_master_address),     //     avalon_master.address
		.master_write            (write_master_avalon_master_write),       //                  .write
		.master_byteenable       (write_master_avalon_master_byteenable),  //                  .byteenable
		.master_writedata        (write_master_avalon_master_writedata),   //                  .writedata
		.master_burstcount       (write_master_avalon_master_burstcount),  //                  .burstcount
		.master_waitrequest      (write_master_avalon_master_waitrequest), //                  .waitrequest
		.control_fixed_location  (write_master_control_fixed_location),    //           control.export
		.control_write_base      (write_master_control_write_base),        //                  .export
		.control_write_length    (write_master_control_write_length),      //                  .export
		.control_go              (write_master_control_go),                //                  .export
		.control_done            (write_master_control_done),              //                  .export
		.user_write_buffer       (write_master_stream_write_buffer),       //              user.export
		.user_buffer_input_data  (write_master_stream_buffer_input_data),  //                  .export
		.user_buffer_full        (write_master_stream_buffer_full),        //                  .export
		.master_read             (),                                       //       (terminated)
		.master_readdata         (16'b0000000000000000),                   //       (terminated)
		.master_readdatavalid    (1'b0),                                   //       (terminated)
		.control_read_base       (32'b00000000000000000000000000000000),   //       (terminated)
		.control_read_length     (32'b00000000000000000000000000000000),   //       (terminated)
		.control_early_done      (),                                       //       (terminated)
		.user_read_buffer        (1'b0),                                   //       (terminated)
		.user_buffer_output_data (),                                       //       (terminated)
		.user_data_available     ()                                        //       (terminated)
	);

	top_LPC_FPGA_mm_interconnect_0 mm_interconnect_0 (
		.clk_divide_8k_0_clock_out_clk                               (clk_divide_8k_0_clock_out_clk),                             //                             clk_divide_8k_0_clock_out.clk
		.DDR3_interface_mp_cmd_reset_n_1_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                            // DDR3_interface_mp_cmd_reset_n_1_reset_bridge_in_reset.reset
		.read_master_clock_reset_reset_reset_bridge_in_reset_reset   (rst_controller_reset_out_reset),                            //   read_master_clock_reset_reset_reset_bridge_in_reset.reset
		.read_master_avalon_master_address                           (read_master_avalon_master_address),                         //                             read_master_avalon_master.address
		.read_master_avalon_master_waitrequest                       (read_master_avalon_master_waitrequest),                     //                                                      .waitrequest
		.read_master_avalon_master_burstcount                        (read_master_avalon_master_burstcount),                      //                                                      .burstcount
		.read_master_avalon_master_byteenable                        (read_master_avalon_master_byteenable),                      //                                                      .byteenable
		.read_master_avalon_master_read                              (read_master_avalon_master_read),                            //                                                      .read
		.read_master_avalon_master_readdata                          (read_master_avalon_master_readdata),                        //                                                      .readdata
		.read_master_avalon_master_readdatavalid                     (read_master_avalon_master_readdatavalid),                   //                                                      .readdatavalid
		.DDR3_interface_avl_1_address                                (mm_interconnect_0_ddr3_interface_avl_1_address),            //                                  DDR3_interface_avl_1.address
		.DDR3_interface_avl_1_write                                  (mm_interconnect_0_ddr3_interface_avl_1_write),              //                                                      .write
		.DDR3_interface_avl_1_read                                   (mm_interconnect_0_ddr3_interface_avl_1_read),               //                                                      .read
		.DDR3_interface_avl_1_readdata                               (mm_interconnect_0_ddr3_interface_avl_1_readdata),           //                                                      .readdata
		.DDR3_interface_avl_1_writedata                              (mm_interconnect_0_ddr3_interface_avl_1_writedata),          //                                                      .writedata
		.DDR3_interface_avl_1_beginbursttransfer                     (mm_interconnect_0_ddr3_interface_avl_1_beginbursttransfer), //                                                      .beginbursttransfer
		.DDR3_interface_avl_1_burstcount                             (mm_interconnect_0_ddr3_interface_avl_1_burstcount),         //                                                      .burstcount
		.DDR3_interface_avl_1_byteenable                             (mm_interconnect_0_ddr3_interface_avl_1_byteenable),         //                                                      .byteenable
		.DDR3_interface_avl_1_readdatavalid                          (mm_interconnect_0_ddr3_interface_avl_1_readdatavalid),      //                                                      .readdatavalid
		.DDR3_interface_avl_1_waitrequest                            (~mm_interconnect_0_ddr3_interface_avl_1_waitrequest)        //                                                      .waitrequest
	);

	top_LPC_FPGA_mm_interconnect_1 mm_interconnect_1 (
		.clk_divide_8k_0_clock_out_clk                               (clk_divide_8k_0_clock_out_clk),                             //                             clk_divide_8k_0_clock_out.clk
		.DDR3_interface_mp_cmd_reset_n_2_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                            // DDR3_interface_mp_cmd_reset_n_2_reset_bridge_in_reset.reset
		.write_master_clock_reset_reset_reset_bridge_in_reset_reset  (rst_controller_reset_out_reset),                            //  write_master_clock_reset_reset_reset_bridge_in_reset.reset
		.write_master_avalon_master_address                          (write_master_avalon_master_address),                        //                            write_master_avalon_master.address
		.write_master_avalon_master_waitrequest                      (write_master_avalon_master_waitrequest),                    //                                                      .waitrequest
		.write_master_avalon_master_burstcount                       (write_master_avalon_master_burstcount),                     //                                                      .burstcount
		.write_master_avalon_master_byteenable                       (write_master_avalon_master_byteenable),                     //                                                      .byteenable
		.write_master_avalon_master_write                            (write_master_avalon_master_write),                          //                                                      .write
		.write_master_avalon_master_writedata                        (write_master_avalon_master_writedata),                      //                                                      .writedata
		.DDR3_interface_avl_2_address                                (mm_interconnect_1_ddr3_interface_avl_2_address),            //                                  DDR3_interface_avl_2.address
		.DDR3_interface_avl_2_write                                  (mm_interconnect_1_ddr3_interface_avl_2_write),              //                                                      .write
		.DDR3_interface_avl_2_read                                   (mm_interconnect_1_ddr3_interface_avl_2_read),               //                                                      .read
		.DDR3_interface_avl_2_readdata                               (mm_interconnect_1_ddr3_interface_avl_2_readdata),           //                                                      .readdata
		.DDR3_interface_avl_2_writedata                              (mm_interconnect_1_ddr3_interface_avl_2_writedata),          //                                                      .writedata
		.DDR3_interface_avl_2_beginbursttransfer                     (mm_interconnect_1_ddr3_interface_avl_2_beginbursttransfer), //                                                      .beginbursttransfer
		.DDR3_interface_avl_2_burstcount                             (mm_interconnect_1_ddr3_interface_avl_2_burstcount),         //                                                      .burstcount
		.DDR3_interface_avl_2_byteenable                             (mm_interconnect_1_ddr3_interface_avl_2_byteenable),         //                                                      .byteenable
		.DDR3_interface_avl_2_readdatavalid                          (mm_interconnect_1_ddr3_interface_avl_2_readdatavalid),      //                                                      .readdatavalid
		.DDR3_interface_avl_2_waitrequest                            (~mm_interconnect_1_ddr3_interface_avl_2_waitrequest)        //                                                      .waitrequest
	);

	top_LPC_FPGA_mm_interconnect_2 mm_interconnect_2 (
		.clk_divide_8k_0_clock_out_clk                             (clk_divide_8k_0_clock_out_clk),                                             //                           clk_divide_8k_0_clock_out.clk
		.avmm_master_interface_0_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                                            // avmm_master_interface_0_reset_reset_bridge_in_reset.reset
		.JTAG_master_clk_reset_reset_bridge_in_reset_reset         (rst_controller_reset_out_reset),                                            //         JTAG_master_clk_reset_reset_bridge_in_reset.reset
		.JTAG_master_master_address                                (jtag_master_master_address),                                                //                                  JTAG_master_master.address
		.JTAG_master_master_waitrequest                            (jtag_master_master_waitrequest),                                            //                                                    .waitrequest
		.JTAG_master_master_byteenable                             (jtag_master_master_byteenable),                                             //                                                    .byteenable
		.JTAG_master_master_read                                   (jtag_master_master_read),                                                   //                                                    .read
		.JTAG_master_master_readdata                               (jtag_master_master_readdata),                                               //                                                    .readdata
		.JTAG_master_master_readdatavalid                          (jtag_master_master_readdatavalid),                                          //                                                    .readdatavalid
		.JTAG_master_master_write                                  (jtag_master_master_write),                                                  //                                                    .write
		.JTAG_master_master_writedata                              (jtag_master_master_writedata),                                              //                                                    .writedata
		.AlgorithmRun_s1_address                                   (mm_interconnect_2_algorithmrun_s1_address),                                 //                                     AlgorithmRun_s1.address
		.AlgorithmRun_s1_write                                     (mm_interconnect_2_algorithmrun_s1_write),                                   //                                                    .write
		.AlgorithmRun_s1_readdata                                  (mm_interconnect_2_algorithmrun_s1_readdata),                                //                                                    .readdata
		.AlgorithmRun_s1_writedata                                 (mm_interconnect_2_algorithmrun_s1_writedata),                               //                                                    .writedata
		.AlgorithmRun_s1_chipselect                                (mm_interconnect_2_algorithmrun_s1_chipselect),                              //                                                    .chipselect
		.avmm_master_interface_0_avmm_master_interface_address     (mm_interconnect_2_avmm_master_interface_0_avmm_master_interface_address),   //       avmm_master_interface_0_avmm_master_interface.address
		.avmm_master_interface_0_avmm_master_interface_write       (mm_interconnect_2_avmm_master_interface_0_avmm_master_interface_write),     //                                                    .write
		.avmm_master_interface_0_avmm_master_interface_read        (mm_interconnect_2_avmm_master_interface_0_avmm_master_interface_read),      //                                                    .read
		.avmm_master_interface_0_avmm_master_interface_readdata    (mm_interconnect_2_avmm_master_interface_0_avmm_master_interface_readdata),  //                                                    .readdata
		.avmm_master_interface_0_avmm_master_interface_writedata   (mm_interconnect_2_avmm_master_interface_0_avmm_master_interface_writedata), //                                                    .writedata
		.DDR3_interface_avl_0_address                              (mm_interconnect_2_ddr3_interface_avl_0_address),                            //                                DDR3_interface_avl_0.address
		.DDR3_interface_avl_0_write                                (mm_interconnect_2_ddr3_interface_avl_0_write),                              //                                                    .write
		.DDR3_interface_avl_0_read                                 (mm_interconnect_2_ddr3_interface_avl_0_read),                               //                                                    .read
		.DDR3_interface_avl_0_readdata                             (mm_interconnect_2_ddr3_interface_avl_0_readdata),                           //                                                    .readdata
		.DDR3_interface_avl_0_writedata                            (mm_interconnect_2_ddr3_interface_avl_0_writedata),                          //                                                    .writedata
		.DDR3_interface_avl_0_beginbursttransfer                   (mm_interconnect_2_ddr3_interface_avl_0_beginbursttransfer),                 //                                                    .beginbursttransfer
		.DDR3_interface_avl_0_burstcount                           (mm_interconnect_2_ddr3_interface_avl_0_burstcount),                         //                                                    .burstcount
		.DDR3_interface_avl_0_byteenable                           (mm_interconnect_2_ddr3_interface_avl_0_byteenable),                         //                                                    .byteenable
		.DDR3_interface_avl_0_readdatavalid                        (mm_interconnect_2_ddr3_interface_avl_0_readdatavalid),                      //                                                    .readdatavalid
		.DDR3_interface_avl_0_waitrequest                          (~mm_interconnect_2_ddr3_interface_avl_0_waitrequest)                        //                                                    .waitrequest
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (jtag_master_master_reset_reset), // reset_in0.reset
		.clk            (clk_divide_8k_0_clock_out_clk),  //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (jtag_master_master_reset_reset),     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
