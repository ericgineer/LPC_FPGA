
module LevinsonDurbinTest (
	clk_clk,
	leds_led);	

	input		clk_clk;
	output	[7:0]	leds_led;
endmodule
